CONFIGURATION WordMux2_untitled_config OF WordMux2 IS
   FOR untitled
   END FOR;
END WordMux2_untitled_config;