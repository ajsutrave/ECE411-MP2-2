ARCHITECTURE UNTITLED OF MEMORY IS
SIGNAL PRE_MEMRESP_H : STD_LOGIC;
SIGNAL PRE_DATAIN : LC3B_WORD;
BEGIN
  -------------------------------------------------------------------
  VHDL_MEMORY : PROCESS (RESET_L, MEMREAD_L, MEMWRITEH_L, MEMWRITEL_L) 
  -------------------------------------------------------------------
  VARIABLE MEM : MEMORY_ARRAY_64K;
  VARIABLE INT_OLD_ADDRESS : INTEGER;
  VARIABLE INT_ADDRESS : INTEGER;
  BEGIN
	  INT_ADDRESS := TO_INTEGER(UNSIGNED('0' & ADDRESS(11 DOWNTO 1) & '0'));
	  IF RESET_L = '0' THEN
		  PRE_MEMRESP_H <= '0';
		  MYDRAMINIT_64K(MEM);
    ELSIF (RESET_L = 'U') AND (MEMREAD_L = 'U') AND (MEMWRITEH_L = 'U') AND (MEMWRITEL_L = 'U') THEN
      -- resetting
      ASSERT TRUE;
	  ELSE
		  IF ((INT_ADDRESS >= 0) AND (INT_ADDRESS <= 4095)) THEN
			  IF (MEMWRITEH_L'EVENT AND (MEMWRITEH_L = '0') AND (MEMWRITEH_L'LAST_VALUE /= '1')) THEN
				  ASSERT FALSE 
				  REPORT "MEMORY WRITE HI-LO TIMING ERROR"
				  SEVERITY FAILURE;
			  END IF;
			  IF (MEMWRITEL_L'EVENT AND (MEMWRITEL_L = '0') AND (MEMWRITEL_L'LAST_VALUE /= '1')) THEN
				  ASSERT FALSE 
				  REPORT "MEMORY WRITE LO-HI TIMING ERROR"
				  SEVERITY FAILURE;
			  END IF;
			  IF (MEMWRITEL_L'EVENT AND (MEMWRITEL_L'LAST_VALUE = '0') AND (INT_ADDRESS /= INT_OLD_ADDRESS)) THEN
				  ASSERT FALSE 
				  REPORT "MEMORY WRITE LO TIMING ERROR"
				  SEVERITY FAILURE;
			  END IF;
			  IF (MEMWRITEH_L'EVENT AND (MEMWRITEH_L'LAST_VALUE = '0') AND (INT_ADDRESS /= INT_OLD_ADDRESS)) THEN
				  ASSERT FALSE 
				  REPORT "MEMORY WRITE HI TIMING ERROR"
				  SEVERITY FAILURE;
			  END IF;
			  IF (MEMREAD_L'EVENT AND (MEMREAD_L'LAST_VALUE = '0') AND (INT_ADDRESS /= INT_OLD_ADDRESS)) THEN
				  ASSERT FALSE 
				  REPORT "MEMORY READ TIMING ERROR"
				  SEVERITY FAILURE;
			  END IF;
			  IF (MEMREAD_L = '0' AND MEMWRITEL_L = '1' AND MEMWRITEH_L = '1') THEN
				  PRE_DATAIN(7 DOWNTO 0) <= MEM(INT_ADDRESS);             
				  PRE_DATAIN(15 DOWNTO 8) <= MEM(INT_ADDRESS + 1);             
				  PRE_MEMRESP_H <= '1' AFTER 0 NS, '0' AFTER CLOCK_PERIOD;
					INT_OLD_ADDRESS := INT_ADDRESS;
			  ELSIF ((MEMWRITEL_L = '0' OR MEMWRITEH_L = '0') AND MEMREAD_L = '1') THEN
				  IF (MEMWRITEL_L = '0') THEN
					  MEM(INT_ADDRESS) := DATAOUT(7 DOWNTO 0);
				  END IF;
				  IF (MEMWRITEH_L = '0') THEN
					  MEM(INT_ADDRESS + 1) := DATAOUT(15 DOWNTO 8);
				  END IF;
				  IF(MEMWRITEH_L = '0' OR MEMWRITEL_L = '0') THEN
					  PRE_MEMRESP_H <= '1' AFTER 0 NS, '0' AFTER CLOCK_PERIOD;
				  END IF;
					INT_OLD_ADDRESS := INT_ADDRESS;
				ELSIF (RESET_L'event AND ((RESET_L = '0') OR (RESET_L = '1'))) THEN
					-- reset_l signal going inactive
					ASSERT TRUE;
				ELSIF (MEMREAD_L'event AND ((MEMREAD_L = '1') AND (MEMREAD_L'LAST_VALUE = '0'))) THEN
					-- read_l signal going inactive
					ASSERT TRUE;
				ELSIF (MEMWRITEL_L'event AND ((MEMWRITEL_L = '1') AND (MEMWRITEL_L'LAST_VALUE = '0'))) THEN
					-- read_l signal going inactive
					ASSERT TRUE;
				ELSIF (MEMWRITEH_L'event AND ((MEMWRITEH_L = '1') AND (MEMWRITEH_L'LAST_VALUE = '0'))) THEN
					-- read_l signal going inactive
					ASSERT TRUE;
				ELSE
				  ASSERT FALSE 
				  REPORT "MEMORY WRITE"
				  SEVERITY FAILURE;
			  END IF;
		  ELSE
			  ASSERT FALSE
			  REPORT "INVALID ADDRESS"
			  SEVERITY FAILURE;
		  END IF;
	  END IF;
  END PROCESS VHDL_MEMORY;
  MEMRESP_H <= PRE_MEMRESP_H'DELAYED(DELAY_MP1_MEM);
  DATAIN <= PRE_DATAIN'DELAYED(DELAY_MP1_MEM);
END ARCHITECTURE untitled;
