CONFIGURATION Reg16_untitled_config OF Reg16 IS
   FOR untitled
   END FOR;
END Reg16_untitled_config;