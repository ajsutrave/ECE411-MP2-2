CONFIGURATION IR_untitled_config OF IR IS
   FOR untitled
   END FOR;
END IR_untitled_config;