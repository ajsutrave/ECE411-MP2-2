CONFIGURATION GenCC_untitled_config OF GenCC IS
   FOR untitled
   END FOR;
END GenCC_untitled_config;