--
-- VHDL Architecture ece411.testblack.untitled
--
-- Created:
--          by - sutrave1.ews (gelib-057-01.ews.illinois.edu)
--          at - 17:27:21 01/24/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
ARCHITECTURE untitled OF testblack IS
BEGIN
END ARCHITECTURE untitled;

